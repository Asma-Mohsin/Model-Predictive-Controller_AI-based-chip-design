VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO traffic_controller
  CLASS BLOCK ;
  FOREIGN traffic_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 280.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END clk
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END enable
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.000 25.200 280.000 25.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.000 74.840 280.000 75.440 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.000 124.480 280.000 125.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.000 174.120 280.000 174.720 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.000 223.760 280.000 224.360 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.000 273.400 280.000 274.000 ;
    END
  END io_oeb[5]
  PIN road1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END road1_out[0]
  PIN road1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END road1_out[1]
  PIN road1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END road1_out[2]
  PIN road2_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END road2_out[0]
  PIN road2_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END road2_out[1]
  PIN road2_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END road2_out[2]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END rst_n
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 274.160 288.405 ;
      LAYER met1 ;
        RECT 4.670 10.640 275.470 288.560 ;
      LAYER met2 ;
        RECT 4.690 10.695 275.450 288.505 ;
      LAYER met3 ;
        RECT 4.000 283.920 276.000 288.485 ;
        RECT 4.400 282.520 276.000 283.920 ;
        RECT 4.000 274.400 276.000 282.520 ;
        RECT 4.000 273.000 275.600 274.400 ;
        RECT 4.000 250.600 276.000 273.000 ;
        RECT 4.400 249.200 276.000 250.600 ;
        RECT 4.000 224.760 276.000 249.200 ;
        RECT 4.000 223.360 275.600 224.760 ;
        RECT 4.000 217.280 276.000 223.360 ;
        RECT 4.400 215.880 276.000 217.280 ;
        RECT 4.000 183.960 276.000 215.880 ;
        RECT 4.400 182.560 276.000 183.960 ;
        RECT 4.000 175.120 276.000 182.560 ;
        RECT 4.000 173.720 275.600 175.120 ;
        RECT 4.000 150.640 276.000 173.720 ;
        RECT 4.400 149.240 276.000 150.640 ;
        RECT 4.000 125.480 276.000 149.240 ;
        RECT 4.000 124.080 275.600 125.480 ;
        RECT 4.000 117.320 276.000 124.080 ;
        RECT 4.400 115.920 276.000 117.320 ;
        RECT 4.000 84.000 276.000 115.920 ;
        RECT 4.400 82.600 276.000 84.000 ;
        RECT 4.000 75.840 276.000 82.600 ;
        RECT 4.000 74.440 275.600 75.840 ;
        RECT 4.000 50.680 276.000 74.440 ;
        RECT 4.400 49.280 276.000 50.680 ;
        RECT 4.000 26.200 276.000 49.280 ;
        RECT 4.000 24.800 275.600 26.200 ;
        RECT 4.000 17.360 276.000 24.800 ;
        RECT 4.400 15.960 276.000 17.360 ;
        RECT 4.000 10.715 276.000 15.960 ;
      LAYER met4 ;
        RECT 10.415 222.535 20.640 284.065 ;
        RECT 23.040 222.535 33.745 284.065 ;
  END
END traffic_controller
END LIBRARY

